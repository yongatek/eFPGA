module mult(aa, bb, out);

input  [17 : 0] aa;
input  [17 : 0] bb;
output [35 : 0] out;

assign out = aa * bb;

endmodule









